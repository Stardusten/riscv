// module alu_ctl(
//     input
// )